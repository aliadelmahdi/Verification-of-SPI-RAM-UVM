
package SPI_test_pkg;

    import uvm_pkg::*;
    import SPI_env_pkg::*;
    import shared_pkg::*;
    import SPI_config_pkg::*;
    import SPI_slave_main_sequence_pkg::*;
    import SPI_ram_sequences_pkg::*;
    import SPI_slave_seq_item_pkg::*;
    import SPI_ram_seq_item_pkg::*;

    `include "SPI_test_base.sv"

    
endpackage : SPI_test_pkg