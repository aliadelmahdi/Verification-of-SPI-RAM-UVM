package SPI_test_pkg;

    import uvm_pkg::*;
    import SPI_env_pkg::*;
    import shared_pkg::*;

    `include "SPI_test_base.sv"

    
endpackage : SPI_test_pkg