`ifndef SPI_SLAVE_PKG_SV
`define SPI_SLAVE_PKG_SV

    `include "SPI_slave_seq_item.sv"
    `include "SPI_slave_sequences.sv"
    `include "SPI_slave_driver.sv"
    `include "SPI_slave_monitor.sv"
    `include "SPI_slave_sequencer.sv"
    `include "SPI_slave_agent.sv"

`endif // SPI_SLAVE_PKG_SV