`ifndef SPI_RAM_SEQUENCES_PKG_SV
`define SPI_RAM_SEQUENCES_PKG_SV

    `include "SPI_ram_main_sequence.sv"
    `include "SPI_ram_reset_sequence.sv"

`endif
