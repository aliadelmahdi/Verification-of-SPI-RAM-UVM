`ifndef SPI_RAM_PKG_SV
`define SPI_RAM_PKG_SV

    `include "SPI_ram_seq_item.sv"
    `include "SPI_ram_sequences.sv"
    `include "SPI_ram_driver.sv"
    `include "SPI_ram_monitor.sv"
    `include "SPI_ram_sequencer.sv"
    `include "SPI_ram_agent.sv"


`endif // SPI_RAM_PKG_SV